module counter();
//complete code
endmodule
