module dotprod();
//complete code
endmodule
