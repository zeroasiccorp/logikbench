module bnand();
//complete code
endmodule
