module addsub();
//complete code
endmodule
