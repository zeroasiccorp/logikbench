module mac();
//complete code
endmodule
