module onehot();
//complete code
endmodule
