module umidev();
//complete code
endmodule
