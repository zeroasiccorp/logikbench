module sum();
//complete code
endmodule
