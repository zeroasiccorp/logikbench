module priority();
//complete code
endmodule
