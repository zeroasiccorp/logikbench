module cordic();
//complete code
endmodule
