module sqdiff();
//complete code
endmodule
