module round();
//complete code
endmodule
