module sqrt();
//complete code
endmodule
