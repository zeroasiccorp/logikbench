module min();
//complete code
endmodule
