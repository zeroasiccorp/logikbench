module sad8x8();
//complete code
endmodule
