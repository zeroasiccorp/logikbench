module fftc();
//complete code
endmodule
