module shifl();
//complete code
endmodule
