module axixbar();
//complete code
endmodule
