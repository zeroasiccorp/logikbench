module abs();
//complete code
endmodule
