module ibex();
//complete code
endmodule
