module absdiff();
//complete code
endmodule
