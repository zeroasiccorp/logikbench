module axihost();
//complete code
endmodule
