module regfile();
//complete code
endmodule
