module rstasync();
//complete code
endmodule
