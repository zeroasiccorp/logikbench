module apbdev();
//complete code
endmodule
