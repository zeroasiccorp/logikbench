module serv();
//complete code
endmodule
