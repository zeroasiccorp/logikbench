module shiftreg ();

// simple shift register

endmodule
