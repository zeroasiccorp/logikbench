module fftr();
//complete code
endmodule
