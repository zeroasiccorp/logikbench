module relu();
//complete code
endmodule
