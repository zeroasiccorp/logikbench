module pipeline();
//complete code
endmodule
