module matmul();
//complete code
endmodule
