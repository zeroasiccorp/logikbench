module crc32();
//complete code
endmodule
