module fifosync();
//complete code
endmodule
