module sobel3x3();
//complete code
endmodule
