module ofdm();
//complete code
endmodule
