module csa();
//complete code
endmodule
