module shiftreg();
//complete code
endmodule
