module umihost();
//complete code
endmodule
