module bxor();
//complete code
endmodule
