module spi();
//complete code
endmodule
