module arbiter();
//complete code
endmodule
