module lfsr();
//complete code
endmodule
