module ialu();
//complete code
endmodule
