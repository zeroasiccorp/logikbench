localparam [8*256-1:0] SINETABLE_256 = {
    8'd125,
    8'd122,
    8'd119,
    8'd116,
    8'd112,
    8'd109,
    8'd106,
    8'd103,
    8'd100,
    8'd97,
    8'd94,
    8'd91,
    8'd88,
    8'd85,
    8'd82,
    8'd79,
    8'd77,
    8'd74,
    8'd71,
    8'd68,
    8'd65,
    8'd63,
    8'd60,
    8'd57,
    8'd55,
    8'd52,
    8'd50,
    8'd47,
    8'd45,
    8'd43,
    8'd40,
    8'd38,
    8'd36,
    8'd34,
    8'd32,
    8'd30,
    8'd28,
    8'd26,
    8'd24,
    8'd22,
    8'd21,
    8'd19,
    8'd17,
    8'd16,
    8'd15,
    8'd13,
    8'd12,
    8'd11,
    8'd10,
    8'd8,
    8'd7,
    8'd6,
    8'd6,
    8'd5,
    8'd4,
    8'd3,
    8'd3,
    8'd2,
    8'd2,
    8'd2,
    8'd1,
    8'd1,
    8'd1,
    8'd1,
    8'd1,
    8'd1,
    8'd1,
    8'd2,
    8'd2,
    8'd2,
    8'd3,
    8'd3,
    8'd4,
    8'd5,
    8'd6,
    8'd6,
    8'd7,
    8'd8,
    8'd10,
    8'd11,
    8'd12,
    8'd13,
    8'd15,
    8'd16,
    8'd17,
    8'd19,
    8'd21,
    8'd22,
    8'd24,
    8'd26,
    8'd28,
    8'd30,
    8'd32,
    8'd34,
    8'd36,
    8'd38,
    8'd40,
    8'd43,
    8'd45,
    8'd47,
    8'd50,
    8'd52,
    8'd55,
    8'd57,
    8'd60,
    8'd63,
    8'd65,
    8'd68,
    8'd71,
    8'd74,
    8'd77,
    8'd79,
    8'd82,
    8'd85,
    8'd88,
    8'd91,
    8'd94,
    8'd97,
    8'd100,
    8'd103,
    8'd106,
    8'd109,
    8'd112,
    8'd116,
    8'd119,
    8'd122,
    8'd125,
    8'd128,
    8'd131,
    8'd134,
    8'd137,
    8'd140,
    8'd144,
    8'd147,
    8'd150,
    8'd153,
    8'd156,
    8'd159,
    8'd162,
    8'd165,
    8'd168,
    8'd171,
    8'd174,
    8'd177,
    8'd179,
    8'd182,
    8'd185,
    8'd188,
    8'd191,
    8'd193,
    8'd196,
    8'd199,
    8'd201,
    8'd204,
    8'd206,
    8'd209,
    8'd211,
    8'd213,
    8'd216,
    8'd218,
    8'd220,
    8'd222,
    8'd224,
    8'd226,
    8'd228,
    8'd230,
    8'd232,
    8'd234,
    8'd235,
    8'd237,
    8'd239,
    8'd240,
    8'd241,
    8'd243,
    8'd244,
    8'd245,
    8'd246,
    8'd248,
    8'd249,
    8'd250,
    8'd250,
    8'd251,
    8'd252,
    8'd253,
    8'd253,
    8'd254,
    8'd254,
    8'd254,
    8'd255,
    8'd255,
    8'd255,
    8'd255,
    8'd255,
    8'd255,
    8'd255,
    8'd254,
    8'd254,
    8'd254,
    8'd253,
    8'd253,
    8'd252,
    8'd251,
    8'd250,
    8'd250,
    8'd249,
    8'd248,
    8'd246,
    8'd245,
    8'd244,
    8'd243,
    8'd241,
    8'd240,
    8'd239,
    8'd237,
    8'd235,
    8'd234,
    8'd232,
    8'd230,
    8'd228,
    8'd226,
    8'd224,
    8'd222,
    8'd220,
    8'd218,
    8'd216,
    8'd213,
    8'd211,
    8'd209,
    8'd206,
    8'd204,
    8'd201,
    8'd199,
    8'd196,
    8'd193,
    8'd191,
    8'd188,
    8'd185,
    8'd182,
    8'd179,
    8'd177,
    8'd174,
    8'd171,
    8'd168,
    8'd165,
    8'd162,
    8'd159,
    8'd156,
    8'd153,
    8'd150,
    8'd147,
    8'd144,
    8'd140,
    8'd137,
    8'd134,
    8'd131,
    8'd128
};
