module gray();
//complete code
endmodule
