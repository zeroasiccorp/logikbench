module rom();
//complete code
endmodule
