module sub();
//complete code
endmodule
