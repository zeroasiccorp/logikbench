module fpu34();
//complete code
endmodule
