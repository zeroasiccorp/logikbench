module fifoasync();
//complete code
endmodule
