/*******************************************************************************
 * Function:  UMI UART Controller
 * Author:    Wenting Zhang
 * Copyright: (c) 2023 Zero ASIC. All rights reserved.
 *
 * License: GNU Lesser General Public License 2.1
 *
 * This module is adapted from the OpenCores UART 16550 compatible controller,
 * the original copyright information is included below.
 ******************************************************************************/

//////////////////////////////////////////////////////////////////////
////                                                              ////
////  uart_rfifo.v (Modified from uart_fifo.v)                    ////
////                                                              ////
////                                                              ////
////  This file is part of the "UART 16550 compatible" project    ////
////  http://www.opencores.org/cores/uart16550/                   ////
////                                                              ////
////  Documentation related to this project:                      ////
////  - http://www.opencores.org/cores/uart16550/                 ////
////                                                              ////
////  Projects compatibility:                                     ////
////  - WISHBONE                                                  ////
////  RS232 Protocol                                              ////
////  16550D uart (mostly supported)                              ////
////                                                              ////
////  Overview (main Features):                                   ////
////  UART core receiver FIFO                                     ////
////                                                              ////
////  To Do:                                                      ////
////  Nothing.                                                    ////
////                                                              ////
////  Author(s):                                                  ////
////      - gorban@opencores.org                                  ////
////      - Jacob Gorban                                          ////
////      - Igor Mohor (igorm@opencores.org)                      ////
////                                                              ////
////  Created:        2001/05/12                                  ////
////  Last Updated:   2002/07/22                                  ////
////                  (See log for the revision history)          ////
////                                                              ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
////                                                              ////
//// Copyright (C) 2000, 2001 Authors                             ////
////                                                              ////
//// This source file may be used and distributed without         ////
//// restriction provided that this copyright statement is not    ////
//// removed from the file and that any derivative work contains  ////
//// the original copyright notice and the associated disclaimer. ////
////                                                              ////
//// This source file is free software; you can redistribute it   ////
//// and/or modify it under the terms of the GNU Lesser General   ////
//// Public License as published by the Free Software Foundation; ////
//// either version 2.1 of the License, or (at your option) any   ////
//// later version.                                               ////
////                                                              ////
//// This source is distributed in the hope that it will be       ////
//// useful, but WITHOUT ANY WARRANTY; without even the implied   ////
//// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ////
//// PURPOSE.  See the GNU Lesser General Public License for more ////
//// details.                                                     ////
////                                                              ////
//// You should have received a copy of the GNU Lesser General    ////
//// Public License along with this source; if not, download it   ////
//// from http://www.opencores.org/lgpl.shtml                     ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
//
// CVS Revision History
//
// $Log: not supported by cvs2svn $
// Revision 1.3  2003/06/11 16:37:47  gorban
// This fixes errors in some cases when data is being read and put to the FIFO at the same time. Patch is submitted by Scott Furman. Update is very recommended.
//
// Revision 1.2  2002/07/29 21:16:18  gorban
// The uart_defines.v file is included again in sources.
//
// Revision 1.1  2002/07/22 23:02:23  gorban
// Bug Fixes:
//  * Possible loss of sync and bad reception of stop bit on slow baud rates fixed.
//   Problem reported by Kenny.Tung.
//  * Bad (or lack of ) loopback handling fixed. Reported by Cherry Withers.
//
// Improvements:
//  * Made FIFO's as general inferable memory where possible.
//  So on FPGA they should be inferred as RAM (Distributed RAM on Xilinx).
//  This saves about 1/3 of the Slice count and reduces P&R and synthesis times.
//
//  * Added optional baudrate output (baud_o).
//  This is identical to BAUDOUT* signal on 16550 chip.
//  It outputs 16xbit_clock_rate - the divided clock.
//  It's disabled by default. Define UART_HAS_BAUDRATE_OUTPUT to use.
//
// Revision 1.16  2001/12/20 13:25:46  mohor
// rx push changed to be only one cycle wide.
//
// Revision 1.15  2001/12/18 09:01:07  mohor
// Bug that was entered in the last update fixed (rx state machine).
//
// Revision 1.14  2001/12/17 14:46:48  mohor
// overrun signal was moved to separate block because many sequential lsr
// reads were preventing data from being written to rx fifo.
// underrun signal was not used and was removed from the project.
//
// Revision 1.13  2001/11/26 21:38:54  gorban
// Lots of fixes:
// Break condition wasn't handled correctly at all.
// LSR bits could lose their values.
// LSR value after reset was wrong.
// Timing of THRE interrupt signal corrected.
// LSR bit 0 timing corrected.
//
// Revision 1.12  2001/11/08 14:54:23  mohor
// Comments in Slovene language deleted, few small fixes for better work of
// old tools. IRQs need to be fix.
//
// Revision 1.11  2001/11/07 17:51:52  gorban
// Heavily rewritten interrupt and LSR subsystems.
// Many bugs hopefully squashed.
//
// Revision 1.10  2001/10/20 09:58:40  gorban
// Small synopsis fixes
//
// Revision 1.9  2001/08/24 21:01:12  mohor
// Things connected to parity changed.
// Clock divider changed.
//
// Revision 1.8  2001/08/24 08:48:10  mohor
// FIFO was not cleared after the data was read bug fixed.
//
// Revision 1.7  2001/08/23 16:05:05  mohor
// Stop bit bug fixed.
// Parity bug fixed.
// WISHBONE read cycle bug fixed,
// OE indicator (Overrun Error) bug fixed.
// PE indicator (Parity Error) bug fixed.
// Register read bug fixed.
//
// Revision 1.3  2001/05/31 20:08:01  gorban
// FIFO changes and other corrections.
//
// Revision 1.3  2001/05/27 17:37:48  gorban
// Fixed many bugs. Updated spec. Changed FIFO files structure. See CHANGES.txt file.
//
// Revision 1.2  2001/05/17 18:34:18  gorban
// First 'stable' release. Should be sythesizable now. Also added new header.
//
// Revision 1.0  2001-05-17 21:27:12+02  jacob
// Initial revision
//
//

`include "uart_defines.vh"

module uart_rfifo #(
    // FIFO parameters
    parameter FIFO_WIDTH = `UART_FIFO_REC_WIDTH,
    parameter FIFO_DEPTH = `UART_FIFO_DEPTH,
    parameter FIFO_POINTER_W = `UART_FIFO_POINTER_W,
    parameter FIFO_COUNTER_W = `UART_FIFO_COUNTER_W
) (
    input clk,
    input nreset,
    input [FIFO_WIDTH-1:0] data_in,
    output [FIFO_WIDTH-1:0] data_out,
    // Control signals
    input push, // push strobe, active high
    input pop, // pop strobe, active high
    // status signals
    output reg overrun,
    output reg [FIFO_COUNTER_W-1:0] count,
    output error_bit,
    input fifo_reset,
    input reset_status
);

    wire [7:0] data8_out;
    // flags FIFO
    reg [2:0] fifo[FIFO_DEPTH-1:0];

    // FIFO pointers
    reg [FIFO_POINTER_W-1:0] top;
    reg [FIFO_POINTER_W-1:0] bottom;

    wire [FIFO_POINTER_W-1:0] top_plus_1 = top + 1'b1;

    uart_raminfr #(FIFO_POINTER_W, 8, FIFO_DEPTH) rfifo (
        .clk (clk),
        .we  (push),
        .a   (top),
        .dpra(bottom),
        .di  (data_in[FIFO_WIDTH-1:FIFO_WIDTH-8]),
        .dpo (data8_out)
    );

    integer i;
    always @(posedge clk or negedge nreset) begin // synchronous FIFO
        if (!nreset) begin
            top <= 0;
            bottom <= 0;
            count <= 0;
            for (i = 0; i < FIFO_DEPTH; i = i + 1) begin
                fifo[i] <= 0;
            end
        end
        else if (fifo_reset) begin
            top <= 0;
            bottom <= 0;
            count <= 0;
            for (i = 0; i < FIFO_DEPTH; i = i + 1) begin
                fifo[i] <= 0;
            end
        end
        else begin
            case ({push, pop})
                2'b10:
                if (count < FIFO_DEPTH)  // overrun condition
                    begin
                    top <= top_plus_1;
                    fifo[top] <= data_in[2:0];
                    count <= count + 1'b1;
                end
                2'b01:
                if (count > 0) begin
                    fifo[bottom] <= 0;
                    bottom <= bottom + 1'b1;
                    count <= count - 1'b1;
                end
                2'b11: begin
                    bottom <= bottom + 1'b1;
                    top <= top_plus_1;
                    fifo[top] <= data_in[2:0];
                end
                default: ;
            endcase
        end
    end  // always

    always @(posedge clk or negedge nreset) begin // synchronous FIFO
        if (!nreset)
            overrun <= 1'b0;
        else if (fifo_reset | reset_status)
            overrun <= 1'b0;
        else if (push & ~pop & (count == FIFO_DEPTH))
            overrun <= 1'b1;
    end  // always


    // please note though that data_out is only valid one clock after pop signal
    assign data_out = {data8_out, fifo[bottom]};

    // Additional logic for detection of error conditions (parity and framing) inside the FIFO
    // for the Line Status Register bit 7
    reg error_det;
    always @(*) begin
        error_det = 1'b0;
        for (i = 0; i < FIFO_DEPTH; i = i + 1) begin
            error_det |= |fifo[i];
        end
    end
    assign error_bit = error_det;

endmodule
