module band();
//complete code
endmodule
