module en8b10b();
//complete code
endmodule
