module l1cache();
//complete code
endmodule
