module viterbi();
//complete code
endmodule
