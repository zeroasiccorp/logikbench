module sine();
//complete code
endmodule
