module median3x3();
//complete code
endmodule
