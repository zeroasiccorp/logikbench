module fpu32();
//complete code
endmodule
