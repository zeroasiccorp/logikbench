module ramdp();
//complete code
endmodule
