module incr();
//complete code
endmodule
