module axidev();
//complete code
endmodule
