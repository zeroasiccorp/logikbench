module rstsync();
//complete code
endmodule
