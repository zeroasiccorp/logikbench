module xbar();
//complete code
endmodule
