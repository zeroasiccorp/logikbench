module rv32dec();
//complete code
endmodule
