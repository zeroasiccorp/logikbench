module ramdist();
//complete code
endmodule
