module shiftb();
//complete code
endmodule
