module mulc();
//complete code
endmodule
