module shiftr();
//complete code
endmodule
