module hamming();
//complete code
endmodule
