module max();
//complete code
endmodule
