module rambm();
//complete code
endmodule
