module bxnor();
//complete code
endmodule
