module conv2d();
//complete code
endmodule
