module cam();
//complete code
endmodule
